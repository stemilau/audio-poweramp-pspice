** Profile: "SCHEMATIC1-freq1"  [ C:\Users\stefa\Desktop\PROIECT1\P1_2022_432A_Stefan_Mihai_AAP_N6_OrCAD\Schematics\proiect-orcad\aap-pspicefiles\schematic1\freq1.sim ] 

** Creating circuit file "freq1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../libraries/1n4148.lib" 
.LIB "../../../libraries/bc817-25.lib" 
.LIB "../../../libraries/bc846b.lib" 
.LIB "../../../libraries/bc856b.lib" 
.LIB "../../../libraries/bzx84c10.lib" 
.LIB "../../../libraries/mjd31cg.lib" 
.LIB "../../../libraries/mjd32cg.lib" 
* From [PSPICE NETLIST] section of C:\Users\stefa\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 0.001ms 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
